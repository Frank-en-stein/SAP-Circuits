CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
11
7 Ground~
168 230 295 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5130 0 0
2
5.89773e-315 0
0
14 Logic Display~
6 186 43 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
391 0 0
2
5.89773e-315 0
0
14 Logic Display~
6 163 45 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
3124 0 0
2
5.89773e-315 0
0
14 Logic Display~
6 140 45 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
3421 0 0
2
5.89773e-315 0
0
14 Logic Display~
6 115 45 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.89773e-315 0
0
14 Logic Display~
6 90 46 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.89773e-315 0
0
14 Logic Display~
6 67 46 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
8901 0 0
2
5.89773e-315 0
0
14 Logic Display~
6 45 47 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
7361 0 0
2
5.89773e-315 0
0
14 Logic Display~
6 22 47 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.89773e-315 0
0
7 74LS173
129 348 102 0 14 29
0 13 4 4 3 7 14 15 8 2
2 16 17 18 19
0
0 0 4832 0
6 74F173
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 512 1 0 0 0
1 U
972 0 0
2
5.89773e-315 0
0
7 74LS173
129 478 109 0 14 29
0 20 4 4 3 5 21 22 6 2
2 23 24 25 26
0
0 0 4832 0
6 74F173
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
5.89773e-315 0
0
14
10 0 2 0 0 4096 0 11 0 0 3 2
516 91
536 91
10 0 2 0 0 4096 0 10 0 0 4 2
386 84
386 267
9 0 2 0 0 0 0 11 0 0 4 4
516 82
536 82
536 254
398 254
9 1 2 0 0 8320 0 10 1 0 0 5
386 75
398 75
398 267
230 267
230 289
4 0 3 0 0 4096 0 11 0 0 7 2
446 109
422 109
0 4 3 0 0 0 0 0 11 7 0 2
440 109
446 109
4 4 3 0 0 12416 0 10 11 0 0 6
316 102
280 102
280 43
415 43
415 109
446 109
2 0 4 0 0 4096 0 11 0 0 10 2
440 91
428 91
2 0 4 0 0 4096 0 10 0 0 10 2
310 84
295 84
3 3 4 0 0 12416 0 10 11 0 0 6
310 93
295 93
295 24
428 24
428 100
440 100
5 1 5 0 0 4224 0 11 2 0 0 3
446 118
186 118
186 61
8 1 6 0 0 4224 0 11 5 0 0 3
446 145
115 145
115 63
5 1 7 0 0 4224 0 10 6 0 0 3
316 111
90 111
90 64
8 1 8 0 0 4224 0 10 9 0 0 3
316 138
22 138
22 65
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
431 12 586 36
436 16 580 32
18 la bar is con here
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
16 389 203 413
21 393 197 409
22 oe1=1 oe2=2 e1=9 e2=10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
229 387 360 411
234 391 354 407
15 d is con to bus
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
382 386 577 410
387 390 571 406
23 d0=14.d1=13.d2=12.d3=11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
18 419 149 443
23 423 143 439
15 q is con to alu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
203 419 366 443
208 423 360 439
19 q0=3 q1=4 q2=5 q3=6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
123 465 278 486
132 472 268 487
17 mr mayb reset pin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
438 35 617 56
447 42 607 57
20 clock pulse con here
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
