CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
5
7 74LS181
132 785 83 0 1 45
0 0
0
0 0 4832 0
7 74LS181
-24 -69 25 -61
2 U3
-7 -70 7 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 0 0 0 0 0
1 U
9172 0 0
2
42655.5 0
0
14 Logic Display~
6 410 819 0 1 2
10 0
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7100 0 0
2
42655.5 0
0
7 74LS173
129 1006 513 0 1 29
0 0
0
0 0 4832 0
6 74F173
-21 -51 21 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 0 0 0 0
1 U
3820 0 0
2
42655.5 0
0
7 74LS173
129 545 514 0 1 29
0 0
0
0 0 4832 0
6 74F173
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 0 0 0 0
1 U
7678 0 0
2
42655.5 0
0
7 74LS157
122 774 331 0 1 29
0 0
0
0 0 4832 0
7 74LS157
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 0 0 0 0
1 U
961 0 0
2
42655.5 0
0
14
10 0 0 0 0 0 0 1 0 0 5 3
747 119
211 119
211 211
12 0 0 0 0 0 0 1 0 0 3 3
747 137
278 137
278 210
11 0 0 0 0 0 0 5 0 0 0 5
806 313
892 313
892 216
278 216
278 207
12 11 0 0 0 0 0 5 1 0 0 6
806 331
821 331
821 263
244 263
244 128
747 128
13 0 0 0 0 0 0 5 0 0 0 5
806 349
837 349
837 230
211 230
211 205
14 9 0 0 0 0 0 5 1 0 0 6
806 367
865 367
865 252
170 252
170 110
747 110
5 2 0 0 0 0 0 3 5 0 0 4
974 522
644 522
644 304
742 304
6 4 0 0 0 0 0 3 5 0 0 4
974 531
676 531
676 322
742 322
7 6 0 0 0 0 0 3 5 0 0 4
974 540
693 540
693 340
742 340
8 8 0 0 0 0 0 3 5 0 0 4
974 549
712 549
712 358
742 358
5 3 0 0 0 0 0 4 5 0 0 4
513 523
423 523
423 313
742 313
6 5 0 0 0 0 0 4 5 0 0 4
513 532
439 532
439 331
742 331
7 7 0 0 0 0 0 4 5 0 0 4
513 541
453 541
453 349
742 349
8 9 0 0 0 0 0 4 5 0 0 4
513 550
472 550
472 367
742 367
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
895 118 1040 139
903 125 1031 140
16 F IS CONN TO BUS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
501 71 686 92
509 78 677 93
21 A IS CONN TO ACCUMLTR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
152 210 185 231
160 217 176 232
2 I3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
196 293 253 314
204 299 244 314
5 W BUS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
921 595 978 616
929 602 969 617
5 C reg
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
584 583 643 604
593 590 633 605
5 B reg
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
